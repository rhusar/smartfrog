<?xml version="1.0"?>
<cdl:cdl xmlns:cdl="http://gridforge.org/cddlm/xml/2004/07/30/"
    xmlns:xs="http://www.w3.org/2001/XMLSchema"
    xmlns:xsi="http://www.w3.org/2001/XMLSchema-instance"
    >
  <cdl:documentation>
    This document declares its elements in the wrong order, so is illegal.
  </cdl:documentation>
    <cdl:system/>
    <cdl:configuration/>
    <cdl:types/>
</cdl:cdl>