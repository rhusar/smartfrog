<?xml version="1.0"?>
<cdl:cdl xmlns:cdl="http://www.gridforum.org/namespaces/2005/02/cddlm/CDL-1.0"
    xmlns:fun="http://smartfrog.org/services/cdl/demo/fun">

  <cdl:import location="classpath:/org/smartfrog/services/cddlm/cdl/demo/fun.cdl"/>


  <cdl:system>

    
    <sound cdl:extends="fun:Sound">
      <filename >c:\music.wav</filename>
      <loops >8</loops>
    </sound>


  </cdl:system>
</cdl:cdl>