<?xml version="1.0"?>
<cdl:cdl xmlns:cdl="http://www.gridforum.org/namespaces/2005/02/cddlm/CDL-1.0"
    xmlns:cmp="http://www.gridforum.org/cddlm/components/2005/02"
    xmlns:sf="http://www.gridforum.org/cddlm/smartfrog/2005/02"
    xmlns:sfi="http://smartfrog.org/types/2006/01/"
    xmlns:base="http://smartfrog.org/services/cdl/base/"
    xmlns:fun="http://smartfrog.org/services/cdl/demo/fun">

  <cdl:import location="classpath:/org/smartfrog/services/cddlm/cdl/cmp/components.cdl"/>

  <!--smartfrog extra classes-->

  <cdl:configuration>

    <!-- Echo something -->
    <fun:Sound cdl:extends="cmp:Component">
      <cmp:CommandPath>org.smartfrog.services.fun.sound.SoundPlayerImpl</cmp:CommandPath>
      <filename sfi:type="trimmed"/>
      <loops sfi:type="integer">1</loops>
      <sfShouldTerminate sfi:type="boolean">true</sfShouldTerminate>
    </fun:Sound>


  </cdl:configuration>
</cdl:cdl>